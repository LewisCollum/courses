package StateBus is
  type StateBus is protected
    
  end type;
end package StateBus;

package body StateBus is
  type StateBus is protected body
                               
                 
  end protected body;
                               
                               
end package StateBus;
