package common is
  type State is (ready, run);
end package;
