library ieee;
use ieee.std_logic_1164;

entity StateController is
  port(
    keypadControl: in KeypadControl
);
end entity StateController;

architecture behavioral of StateController is

end architecture behavioral;
