port(
  control: in I2CControlBus;
  )





process
  control.rw
    control.enable
