library ieee;
use ieee.numeric_std.unsigned;

package DataBus is
  subtype word is unsigned(7 downto 0);
end package;
